module mux16to1(in,sel,out);
  input [15:0]in;
  input [3:0]sel;
  output out;
  wire [3:0]t;

  mux4to1 M0 (in[3:0],sel[1:0],t[0]);
  mux4to1 M0 (in[7:4],sel[1:0],t[1]);
  mux4to1 M0 (in[11:8],sel[1:0],t[2]);
  mux4to1 M0 (in[15:12],sel[1:0],t[3]);
  mux4to1 M5 (t,sel[3:2],out);
endmodule

module mux4to1(in,sel,out);
  input [3:0]in;
  input [1:0]sel;
  ouput out;
  wire [1:0]t;

  mux2to1 M0 (in[1:0],sel[0],t[0]);
  mux2to1 M0 (in[3:2],sel[0],t[1]);
  mux2to1 M0 (t,sel[1],out);
endmodule

module mux2to1 (in,sel,out);
  input [1:0]in;
  input sel;
  output out;
  assign out = in[sel];
endmodule
  
